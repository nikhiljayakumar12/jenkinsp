module design_hello (
input a,
output b
);

assign b=a;
endmodule
